module sap ();
