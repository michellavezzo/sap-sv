//module sap ();